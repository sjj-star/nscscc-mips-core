`define PC_INITIAL 32'hbfc0_0000
`define PC_EBASE   32'hbfc0_0380
`define INST_INTI  32'h0000_0000

`define ADDR_SEG3 3'b111
`define ADDR_SSEG 3'b110
`define ADDR_SEG1 3'b101
`define ADDR_SEG0 3'b100

`define INT 5'h00
`define ADEL 5'h04
`define ADES 5'h05
`define SYS 5'h08
`define BP 5'h09
`define RI 5'h0a
`define OV 5'h0c
`define INVALID_EXCEP 5'h15

//`default_nettype none
