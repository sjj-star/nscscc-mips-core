`undef PC_INITIAL
`undef PC_EBASE
`undef INST_INTI

`undef ADDR_SEG3
`undef ADDR_SSEG
`undef ADDR_SEG1
`undef ADDR_SEG0

`undef INT
`undef ADEL
`undef ADES
`undef SYS
`undef BP
`undef RI
`undef OV
`undef INVALID_EXCEP

//`default_nettype none
